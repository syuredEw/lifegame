module lifegame_cal(
    input       clk, 
    input       rst, 

    input [8:0] neibor,
    input       cal_enable,
    output     outdata
);

    
    logic data;
    assign outdata = data   ;
    always @(posedge clk)
    begin
        if(cal_enable)
        begin
            case( neibor )
                9'b000_000_111: data <= 1'b1;
                9'b000_001_011: data <= 1'b1;
                9'b000_001_101: data <= 1'b1;
                9'b000_001_110: data <= 1'b1;
                9'b000_010_011: data <= 1'b1;
                9'b000_010_101: data <= 1'b1;
                9'b000_010_110: data <= 1'b1;
                9'b000_010_111: data <= 1'b1;
                9'b000_011_001: data <= 1'b1;
                9'b000_011_010: data <= 1'b1;
                9'b000_011_011: data <= 1'b1;
                9'b000_011_100: data <= 1'b1;
                9'b000_011_101: data <= 1'b1;
                9'b000_011_110: data <= 1'b1;
                9'b000_100_011: data <= 1'b1;
                9'b000_100_101: data <= 1'b1;
                9'b000_100_110: data <= 1'b1;
                9'b000_101_001: data <= 1'b1;
                9'b000_101_010: data <= 1'b1;
                9'b000_101_100: data <= 1'b1;
                9'b000_110_001: data <= 1'b1;
                9'b000_110_010: data <= 1'b1;
                9'b000_110_011: data <= 1'b1;
                9'b000_110_100: data <= 1'b1;
                9'b000_110_011: data <= 1'b1;
                9'b000_110_100: data <= 1'b1;
                9'b000_110_101: data <= 1'b1;
                9'b000_110_110: data <= 1'b1;
                9'b000_111_000: data <= 1'b1;
                9'b000_111_001: data <= 1'b1;
                9'b000_111_010: data <= 1'b1;
                9'b000_111_100: data <= 1'b1;
                9'b001_000_101: data <= 1'b1;
                9'b001_000_110: data <= 1'b1;
                9'b001_001_001: data <= 1'b1;
                9'b001_001_010: data <= 1'b1;
                9'b001_001_100: data <= 1'b1;
                9'b001_010_001: data <= 1'b1;
                9'b001_010_010: data <= 1'b1;
                9'b001_010_011: data <= 1'b1;
                9'b001_010_100: data <= 1'b1;
                9'b001_010_101: data <= 1'b1;
                9'b001_010_110: data <= 1'b1;
                9'b001_011_000: data <= 1'b1;
                9'b001_011_001: data <= 1'b1;
                9'b001_011_010: data <= 1'b1;
                9'b001_011_100: data <= 1'b1;
                9'b001_100_001: data <= 1'b1;
                9'b001_100_010: data <= 1'b1;
                9'b001_100_100: data <= 1'b1;
                9'b001_101_000: data <= 1'b1;
                9'b001_110_000: data <= 1'b1;
                9'b001_110_001: data <= 1'b1;
                9'b001_110_010: data <= 1'b1;
                9'b001_110_100: data <= 1'b1;
                9'b001_110_100: data <= 1'b1;
                9'b001_111_000: data <= 1'b1;
                9'b010_000_011: data <= 1'b1;
                9'b010_000_101: data <= 1'b1;
                9'b010_000_110: data <= 1'b1;
                9'b010_001_001: data <= 1'b1;
                9'b010_001_010: data <= 1'b1;
                9'b010_001_100: data <= 1'b1;
                9'b010_010_001: data <= 1'b1;
                9'b010_010_010: data <= 1'b1;
                9'b010_010_011: data <= 1'b1;
                9'b010_010_100: data <= 1'b1;
                9'b010_010_101: data <= 1'b1;
                9'b010_010_110: data <= 1'b1;
                9'b010_011_000: data <= 1'b1;
                9'b010_011_001: data <= 1'b1;
                9'b010_011_010: data <= 1'b1;
                9'b010_011_100: data <= 1'b1;
                9'b010_100_001: data <= 1'b1;
                9'b010_100_010: data <= 1'b1;
                9'b010_100_100: data <= 1'b1;
                9'b010_101_000: data <= 1'b1;
                9'b010_110_000: data <= 1'b1;
                9'b010_110_001: data <= 1'b1;
                9'b010_110_100: data <= 1'b1;
                9'b010_111_000: data <= 1'b1;
                9'b011_000_001: data <= 1'b1;
                9'b011_000_010: data <= 1'b1;
                9'b011_000_100: data <= 1'b1;
                9'b011_001_000: data <= 1'b1;
                9'b011_010_001: data <= 1'b1;
                9'b011_010_001: data <= 1'b1;
                9'b011_010_010: data <= 1'b1;
                9'b011_010_100: data <= 1'b1;
                9'b011_011_000: data <= 1'b1;
                9'b011_100_000: data <= 1'b1;
                9'b011_110_000: data <= 1'b1;
                9'b100_000_011: data <= 1'b1;
                9'b100_000_101: data <= 1'b1;
                9'b100_000_110: data <= 1'b1;
                9'b100_001_001: data <= 1'b1;
                9'b100_001_010: data <= 1'b1;
                9'b100_001_100: data <= 1'b1;
                9'b100_010_001: data <= 1'b1;
                9'b100_010_010: data <= 1'b1;
                9'b100_010_011: data <= 1'b1;
                9'b100_010_100: data <= 1'b1;
                9'b100_010_101: data <= 1'b1;
                9'b100_010_110: data <= 1'b1;
                9'b100_011_000: data <= 1'b1;
                9'b100_011_001: data <= 1'b1;
                9'b100_011_010: data <= 1'b1;
                9'b100_011_100: data <= 1'b1;
                9'b100_100_001: data <= 1'b1;
                9'b100_100_010: data <= 1'b1;
                9'b100_100_100: data <= 1'b1;
                9'b100_110_000: data <= 1'b1;
                9'b100_110_001: data <= 1'b1;
                9'b100_110_010: data <= 1'b1;
                9'b100_110_011: data <= 1'b1;
                9'b100_110_100: data <= 1'b1;
                9'b101_000_001: data <= 1'b1;
                9'b101_000_010: data <= 1'b1;
                9'b101_000_100: data <= 1'b1;
                9'b101_001_000: data <= 1'b1;
                9'b101_010_000: data <= 1'b1;
                9'b101_010_001: data <= 1'b1;
                9'b101_010_010: data <= 1'b1;
                9'b101_010_100: data <= 1'b1;
                9'b101_011_000: data <= 1'b1;
                9'b101_100_000: data <= 1'b1;
                9'b101_110_000: data <= 1'b1;
                9'b110_000_001: data <= 1'b1;
                9'b110_000_010: data <= 1'b1;
                9'b110_000_100: data <= 1'b1;
                9'b110_001_000: data <= 1'b1;
                9'b110_010_000: data <= 1'b1;
                9'b110_010_001: data <= 1'b1;
                9'b110_010_010: data <= 1'b1;
                9'b110_010_100: data <= 1'b1;
                9'b110_011_000: data <= 1'b1;
                9'b110_100_000: data <= 1'b1;
                9'b110_110_000: data <= 1'b1;
                9'b111_000_000: data <= 1'b1;
                9'b110_011_000: data <= 1'b1;
                9'b111_010_000: data <= 1'b1;
                
                default : data <= 1'b0;
            endcase
        end
    end
    
    
endmodule
